-- A DUT entity is used to wrap your design.
--  This example shows how you can do this for the
--  Full-adder.

library ieee;
use ieee.std_logic_1164.all;

entity DUT is
   port(input_vector: in std_logic_vector(5 downto 0);
       	output_vector: out std_logic_vector(0 downto 0));
end entity;

architecture DutWrap of DUT is
	-- Instantiate your own top Module component in place of ALU_1
	Component divisibility is
		port(
				F: in std_logic;
				X: in std_logic_vector(4 downto 0);
			   Y  : out std_logic
			);
	end component divisibility;
begin

   -- input/output vector element ordering is critical,
   -- and must match the ordering in the trace file!
   add_instance: divisibility 
	port map (
	F => input_vector(5), 
	X => input_vector(4 downto 0),
	Y => output_vector(0)
	);

end DutWrap;

